library verilog;
use verilog.vl_types.all;
entity musa is
end musa;
