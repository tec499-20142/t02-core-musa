module musa();


endmodule