module stack ();

endmodule