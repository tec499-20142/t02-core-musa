module ula(
	input [31:0] inA;
	input [31:0] inB;
	input op;
	input fx;
	output [32:0]result;
	output wire overF;
	output wire zero;
);
	

endmodule