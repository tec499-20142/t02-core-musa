module musa();


endmodule